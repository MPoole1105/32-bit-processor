----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Matthew Poole
-- 
-- Create Date: 14.10.2024 17:03:05
-- Design Name: 
-- Module Name: RF_Mux_32_1Bit_2337347_t B- Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity RF_32_1Bit_2337347_TB is
--  Port ( );
end RF_32_1Bit_2337347_TB;

architecture Simulation of RF_Mux_32_1Bit_2337347_TB is
    component RF_Mux_32_1Bit_23373470 
    Port(I0 : in std_logic;  
     I1 : in std_logic;  
     I2 : in std_logic;  
     I3 : in std_logic;  
     I4 : in std_logic;  
     I5 : in std_logic;  
     I6 : in std_logic;  
     I7 : in std_logic;  
     I8 : in std_logic;  
     I9 : in std_logic;  
     I10 : in std_logic; 
     I11 : in std_logic; 
     I12 : in std_logic; 
     I13 : in std_logic; 
     I14 : in std_logic; 
     I15 : in std_logic; 
     I16 : in std_logic; 
     I17 : in std_logic; 
     I18 : in std_logic; 
     I19 : in std_logic; 
     I20 : in std_logic; 
     I21 : in std_logic; 
     I22 : in std_logic; 
     I23 : in std_logic; 
     I24 : in std_logic; 
     I25 : in std_logic; 
     I26 : in std_logic; 
     I27 : in std_logic; 
     I28 : in std_logic; 
     I29 : in std_logic; 
     I30 : in std_logic; 
     I31 : in std_logic; 
     S : in std_logic_vector (4 downto 0);
     Y : out std_logic );
    end component;
        
signal I : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000";  
signal Y_TB : std_logic := '0';
signal S_TB : std_logic_vector (4 downto 0) := b"00000";

constant STUDENTID : std_logic_vector (31 downto 0) := x"0164A69E";

begin
-- Instantiate the Mux
    uut: RF_Mux_32_1Bit_23373470
        Port map (I0 => I(0),
                  I1 => I(1),
                  I2 => I(2),
                  I3 => I(3),
                  I4 => I(4),
                  I5 => I(5),
                  I6 => I(6),
                  I7 => I(7),
                  I8 => I(8),
                  I9 => I(9),
                  I10 => I(10),
                  I11 => I(11),
                  I12 => I(12),
                  I13 => I(13),
                  I14 => I(14),
                  I15 => I(15),
                  I16 => I(16),
                  I17 => I(17),
                  I18 => I(18),
                  I19 => I(19),
                  I20 => I(20),
                  I21 => I(21),
                  I22 => I(22),
                  I23 => I(23),
                  I24 => I(24),
                  I25 => I(25),
                  I26 => I(26),
                  I27 => I(27),
                  I28 => I(28),
                  I29 => I(29),
                  I30 => I(30),
                  I31 => I(31),
                  S => S_TB,
                  Y => Y_TB);
                  
stim_proc: process
   begin		
      S_TB <= "00000";                                            -- case A   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      
      
      wait for 60 ns;
      I(0) <= '1'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "00001";                                            -- case B   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '1'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "00010";                                            -- case C   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '1'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;

      S_TB <= "00011";                                            -- case D   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '1';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;

      S_TB <= "00100";                                            -- case E   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '1'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "00101";                                            -- case F   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '1'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "00110";                                            -- case G   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '1'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;

      S_TB <= "00111";                                            -- case H   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '1';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "01000";                                            -- case A   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      
      
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '1'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "01001";                                            -- case B   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '1'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "01010";                                            -- case C   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '1'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;

      S_TB <= "01011";                                            -- case D   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '1'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;

      S_TB <= "01100";                                            -- case E   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '1'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "01101";                                            -- case F   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '1'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "01110";                                            -- case G   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '1'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;

      S_TB <= "01111";                                            -- case H   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '1'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "10000";                                            -- case A   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      
      
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '1'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "10001";                                            -- case B   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '1'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "10010";                                            -- case C   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '1'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;

      S_TB <= "10011";                                            -- case D   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '1'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;

      S_TB <= "10100";                                            -- case E   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '1'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "10101";                                            -- case F   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '1'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "10110";                                            -- case G   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '1'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;

      S_TB <= "10111";                                            -- case H   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '1';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "11000";                                            -- case A   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      
      
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '1'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "11001";                                            -- case B   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '1'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "11010";                                            -- case C   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '1'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;

      S_TB <= "11011";                                            -- case D   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '1';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;

      S_TB <= "11100";                                            -- case E   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '1'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "11101";                                            -- case F   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '1'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      
      S_TB <= "11110";                                            -- case G   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '1'; I(31) <= '0'; 
      wait for 60 ns;

      S_TB <= "11111";                                            -- case H   
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '0'; 
      wait for 60 ns;
      I(0) <= '0'; I(1) <= '0'; I(2) <= '0'; I(3) <= '0';
      I(4) <= '0'; I(5) <= '0'; I(6) <= '0'; I(7) <= '0';
      I(8) <= '0'; I(9) <= '0'; I(10) <= '0'; I(11) <= '0'; 
      I(12) <= '0'; I(13) <= '0'; I(14) <= '0'; I(15) <= '0'; 
      I(16) <= '0'; I(17) <= '0'; I(18) <= '0'; I(19) <= '0'; 
      I(20) <= '0'; I(21) <= '0'; I(22) <= '0'; I(23) <= '0';
      I(24) <= '0'; I(25) <= '0'; I(26) <= '0'; I(27) <= '0';
      I(28) <= '0'; I(29) <= '0'; I(30) <= '0'; I(31) <= '1'; 
      wait for 60 ns;
      
   end process;


end Simulation;

begin


end Simulation;


-- Company: 
-- Engineer: Matthew Poole
-- 
-- Create Date: 15.10.2024 14:19:48
-- Design Name: 
-- Module Name: RF_Mux_32_32Bit_23373470_TB - Simulation
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity RF_Mux_32_32Bit_23373470_TB is
--  Port ( );
end RF_Mux_32_32Bit_23373470_TB;

architecture Simulation of RF_Mux_32_32Bit_23373470_TB is
component RF_Mux_32_32Bit_23373470 is
Port(I0 : in std_logic_vector (31 downto 0);
         I1 : in std_logic_vector (31 downto 0);
         I2 : in std_logic_vector (31 downto 0);
         I3 : in std_logic_vector (31 downto 0);
         I4 : in std_logic_vector (31 downto 0);
         I5 : in std_logic_vector (31 downto 0);
         I6 : in std_logic_vector (31 downto 0);
         I7 : in std_logic_vector (31 downto 0);
         I8 : in std_logic_vector (31 downto 0);
         I9 : in std_logic_vector (31 downto 0);
         I10 : in std_logic_vector (31 downto 0);
         I11 : in std_logic_vector (31 downto 0);
         I12 : in std_logic_vector (31 downto 0);
         I13 : in std_logic_vector (31 downto 0);
         I14 : in std_logic_vector (31 downto 0);
         I15 : in std_logic_vector (31 downto 0);
         I16 : in std_logic_vector (31 downto 0);
         I17 : in std_logic_vector (31 downto 0);
         I18 : in std_logic_vector (31 downto 0);
         I19 : in std_logic_vector (31 downto 0);
         I20 : in std_logic_vector (31 downto 0);
         I21 : in std_logic_vector (31 downto 0);
         I22 : in std_logic_vector (31 downto 0);
         I23 : in std_logic_vector (31 downto 0);
         I24 : in std_logic_vector (31 downto 0);
         I25 : in std_logic_vector (31 downto 0);
         I26 : in std_logic_vector (31 downto 0);
         I27 : in std_logic_vector (31 downto 0);
         I28 : in std_logic_vector (31 downto 0);
         I29 : in std_logic_vector (31 downto 0);
         I30 : in std_logic_vector (31 downto 0);
         I31 : in std_logic_vector (31 downto 0);
         S : in std_logic_vector (4 downto 0);
         Y : out std_logic_vector (31 downto 0));
         
         
end component;
 signal I0 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I1 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I2 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I3 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000";
 signal I4 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I5 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I6 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I7 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I8 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I9 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I10 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I11 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I12 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I13 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I14 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I15 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I16 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I17 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I18 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I19 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I20 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I21 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I22 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I23 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I24 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I25 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I26 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I27 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I28 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I29 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I30 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 signal I31 : std_logic_vector (31 downto 0) := b"00000000000000000000000000000000"; 
 
 signal S_TB : std_logic_vector (4 downto 0) := b"00000";
 signal Y_TB : std_logic_vector (31 downto 0);
 constant StudentID : STD_LOGIC_VECTOR (27 downto 0) := x"164A69E";  


begin
uut: RF_Mux_32_32Bit_23373470
        Port map (I0 => I0,
                  I1 => I1,
                  I2 => I2,
                  I3 => I3,
                  I4 => I4,
                  I5 => I5,
                  I6 => I6,
                  I7 => I7,
                  I8 => I8,
                  I9 => I9,
                  I10 => I10,
                  I11 => I11,
                  I12 => I12,
                  I13 => I13,
                  I14 => I14,
                  I15 => I15,
                  I16 => I16,
                  I17 => I17,
                  I18 => I18,
                  I19 => I19,
                  I20 => I20,
                  I21 => I21,
                  I22 => I22,
                  I23 => I23,
                  I24 => I24,
                  I25 => I25,
                  I26 => I26,
                  I27 => I27,
                  I28 => I28,
                  I29 => I29,
                  I30 => I30,
                  I31 => I31,
                  S => S_TB,
                  Y => Y_TB);


stim_proc: process
   begin		
      S_TB <= "00000";                                            -- case A   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      
      
      wait for 100 ns;
      I0 <= x"0164A69E"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "00001";                                            -- case B   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= x"0164A69E"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "00010";                                            -- case C   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= x"0164A69E"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;

      S_TB <= "00011";                                            -- case D   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= x"0164A69E";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;

      S_TB <= "00100";                                            -- case E   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= x"0164A69E"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "00101";                                            -- case F   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= x"0164A69E"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "00110";                                            -- case G   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= x"0164A69E"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;

      S_TB <= "00111";                                            -- case H   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= x"0164A69E";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "01000";                                            -- case A   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      
      
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= x"0164A69E"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "01001";                                            -- case B   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= x"0164A69E"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "01010";                                            -- case C   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= x"0164A69E"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;

      S_TB <= "01011";                                            -- case D   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= x"0164A69E"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;

      S_TB <= "01100";                                            -- case E   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= x"0164A69E"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "01101";                                            -- case F   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= x"0164A69E"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "01110";                                            -- case G   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= x"0164A69E"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;

      S_TB <= "01111";                                            -- case H   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= x"0164A69E"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "10000";                                            -- case A   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      
      
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= x"0164A69E"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "10001";                                            -- case B   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= x"0164A69E"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "10010";                                            -- case C   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= x"0164A69E"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;

      S_TB <= "10011";                                            -- case D   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= x"0164A69E"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;

      S_TB <= "10100";                                            -- case E   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= x"0164A69E"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "10101";                                            -- case F   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= x"0164A69E"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "10110";                                            -- case G   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= x"0164A69E"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;

      S_TB <= "10111";                                            -- case H   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= x"0164A69E";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "11000";                                            -- case A   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      
      
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= x"0164A69E"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "11001";                                            -- case B   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= x"0164A69E"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "11010";                                            -- case C   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= x"0164A69E"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;

      S_TB <= "11011";                                            -- case D   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= x"0164A69E";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;

      S_TB <= "11100";                                            -- case E   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= x"0164A69E"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "11101";                                            -- case F   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= x"0164A69E"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      
      S_TB <= "11110";                                            -- case G   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= x"0164A69E"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;

      S_TB <= "11111";                                            -- case H   
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= "00000000000000000000000000000000"; 
      wait for 100 ns;
      I0 <= "00000000000000000000000000000000"; I1 <= "00000000000000000000000000000000"; I2 <= "00000000000000000000000000000000"; I3 <= "00000000000000000000000000000000";
      I4 <= "00000000000000000000000000000000"; I5 <= "00000000000000000000000000000000"; I6 <= "00000000000000000000000000000000"; I7 <= "00000000000000000000000000000000";
      I8 <= "00000000000000000000000000000000"; I9 <= "00000000000000000000000000000000"; I10 <= "00000000000000000000000000000000"; I11 <= "00000000000000000000000000000000"; 
      I12 <= "00000000000000000000000000000000"; I13 <= "00000000000000000000000000000000"; I14 <= "00000000000000000000000000000000"; I15 <= "00000000000000000000000000000000"; 
      I16 <= "00000000000000000000000000000000"; I17 <= "00000000000000000000000000000000"; I18 <= "00000000000000000000000000000000"; I19 <= "00000000000000000000000000000000"; 
      I20 <= "00000000000000000000000000000000"; I21 <= "00000000000000000000000000000000"; I22 <= "00000000000000000000000000000000"; I23 <= "00000000000000000000000000000000";
      I24 <= "00000000000000000000000000000000"; I25 <= "00000000000000000000000000000000"; I26 <= "00000000000000000000000000000000"; I27 <= "00000000000000000000000000000000";
      I28 <= "00000000000000000000000000000000"; I29 <= "00000000000000000000000000000000"; I30 <= "00000000000000000000000000000000"; I31 <= x"0164A69E"; 
      wait for 100 ns;
      
      

   end process;

end Simulation;
